library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity incrementer is
    port (
        clk, rst, en : in std_logic;

    );
end incrementer;

architecture incr of incrementer is
begin

end incr;