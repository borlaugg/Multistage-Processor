library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.basic.all;

entity datapath is
    port (
        
    );
end datapath;

architecture datapath_arch of datapath is

begin

end architecture;